module g3

pub struct Vector2d{
	pub mut:
	x f64
	y f64
	z f64
}
