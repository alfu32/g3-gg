module g3


fn test_entity_interface_casting(){
	entity_interface_casting()
}
fn test_entity_init() {
	entity_init()
}

