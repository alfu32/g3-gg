module main

fn main() {
	v:=[f64(10),10,20,30,40]
	println('Hello World!')
}
